/**********************************************************************************************
 * Project Name       : PISO MODULE
 * Engineer           : Daniel Diaz Platon
 * Module description : An RTL modelling for the transmitter's frame generator,
 *                      and shift register to send data serially in 11 baud_clk cycles.
 * Target             : 5CSXFC6D6F31C6
 * Date               : 2024/05/08
 **********************************************************************************************/

module PISO(
    input wire           reset_n,            //  Active low reset.
    input wire           send,               //  An enable to start sending data.
    input wire           baud_clk,           //  Clocking signal from the BaudGen unit.
    input wire           parity_bit,         //  The parity bit from the Parity unit.
    input wire [1:0]     parity_type,        //  Parity type agreed upon by the Tx and Rx units.
    input wire [7:0]     data_in,            //  The data input.
  
    output reg 	         data_tx, 	         //  Serial transmitter's data out
	output reg 	         active_flag,        //  high when Tx is transmitting, low when idle.
	output reg  	     done_flag 	         //  high when transmission is done, low when active.
);

//  Internal declarations
reg [3:0]   stop_count;
//  an index for the bit of the frame which its turn to get transmitted.
reg [10:0]  frame;
reg [10:0]  frame_r;
//  Holds the data untill transmission is done.
reg         next_state;
//  Holds the FSM's next state.

//  Encoding the states
localparam IDLE   = 1'b0,
           ACTIVE = 1'b1;

//  Frame generation combinational logic
always @(parity_type, parity_bit, data_in)
begin
    if ((~|parity_type) || (&parity_type))
    //  This is an equivalent condition to (parity_type == 'b00)
    //  or (parity_type == 'b11), in order to avoid comparators/xors
    begin
        //  Frame: {idle 1 if needed,stopbit,ParityBit,RegOut[MSB:LSB],Startbit}
        //  Frame with no parity bit
        frame  = {2'b11,data_in,1'b0};
    end
    else
    begin
        //  Frame: {idle 1 if needed,stopbit,ParityBit,RegOut[MSB:LSB],Startbit}
        //  Frame with parity bit
        frame  = {1'b1,parity_bit,data_in,1'b0};
    end
end

//  Transmission logic FSM with Asynchronous Reset logic
always @(posedge baud_clk, negedge reset_n)
begin
    if (~reset_n) 
    begin
       //  idle
        next_state       <= IDLE; 
    end
	else
	begin
		frame_r <= frame;
		case (next_state)

            //  waits for the send enable signal
            IDLE:
            begin
                data_tx      <= 1'b1;
                active_flag  <= 1'b0;
                done_flag    <= 1'b1;
                stop_count   <= 4'd0;

                if (send)
                //  Works as an enable
                begin
                    next_state   <= ACTIVE;
                end
                else
                begin
                    next_state   <= IDLE;
                end
            end

            //  loops 11 time at baud_clk to send all the frame serially
            ACTIVE:
            begin
                if (stop_count[3] && stop_count[1] && stop_count[0])
                //  This is an equivalent condition to (stop_count == 'd11)
                //  in order to avoid comparators/xors  
                begin
                    data_tx      <= 1'b1;
                    stop_count   <= 4'd0;
                    active_flag  <= 1'b0;
                    done_flag    <= 1'b1;
                    next_state   <= IDLE;
                end
                else
                begin
                    data_tx      <= frame_r[0];
                    frame_r      <= frame_r >> 1;
                    //  assiginning the first bit of the frame to the data_tx,
                    //  truncates the rest, then shifting the frame by 1 position
                    //  to the right to get the next data bit, and so on.
                    stop_count   <= stop_count + 1'd1;
                    active_flag  <= 1'b1;
                    done_flag    <= 1'b0;
                    next_state   <= ACTIVE;
                end
            end

            //  Automatically directs to the IDLE state
            default:
            begin
                next_state   <= IDLE;
            end
        endcase 
	end 
end
endmodule  